module EEPROM(
	input	[6:0] Address,	

	
	output reg [17:0]	EEPROM_OUT
);



	always @(*) begin
		case (Address)
			7'bxxxx000: EEPROM_OUT = 18'b000110000000000000;
			7'bxxxx001: EEPROM_OUT = 18'b010000110000000000;
			7'b0000010: EEPROM_OUT = 18'b000000000000000000;
			7'b0000011: EEPROM_OUT = 18'b000000000000000000;
			7'b0000100: EEPROM_OUT = 18'b000000000000000000;
			7'b0001010: EEPROM_OUT = 18'b000010001000000000;
			7'b0001011: EEPROM_OUT = 18'b000000100010000000;
			7'b0001100: EEPROM_OUT = 18'b000000000000000000;
			7'b0010010: EEPROM_OUT = 18'b000000001010000000;
			7'b0010011: EEPROM_OUT = 18'b000000000000000000;
			7'b0010100: EEPROM_OUT = 18'b000000000000000000;
			7'b0011010: EEPROM_OUT = 18'b000010001000000000;
			7'b0011011: EEPROM_OUT = 18'b000001000100000000;
			7'b0011100: EEPROM_OUT = 18'b000000000000000000;
			7'b0100010: EEPROM_OUT = 18'b000010001000000000;
			7'b0100011: EEPROM_OUT = 18'b000000100000000010;
			7'b0100100: EEPROM_OUT = 18'b000000000010001000;
			7'b0101010: EEPROM_OUT = 18'b000010001000000000;
			7'b0101011: EEPROM_OUT = 18'b000000100000000010;
			7'b0101100: EEPROM_OUT = 18'b000000000011001000;
			7'b0110010: EEPROM_OUT = 18'b000010001000000000;
			7'b0110011: EEPROM_OUT = 18'b000000100000000010;
			7'b0110100: EEPROM_OUT = 18'b000000000010011000;
			7'b0111010: EEPROM_OUT = 18'b000010001000000000;
			7'b0111011: EEPROM_OUT = 18'b000000100000000010;
			7'b0111100: EEPROM_OUT = 18'b000000000010101000;
			7'b1000010: EEPROM_OUT = 18'b000010001000000000;
			7'b1000011: EEPROM_OUT = 18'b000000100000000010;
			7'b1000100: EEPROM_OUT = 18'b000000000010111000;
			7'b1001010: EEPROM_OUT = 18'b000000000010111100;
			7'b1001011: EEPROM_OUT = 18'b000000000000000000;
			7'b1001100: EEPROM_OUT = 18'b000000000000000000;
			7'b1010010: EEPROM_OUT = 18'b001000001000000000;
			7'b1010011: EEPROM_OUT = 18'b000000000000000000;
			7'b1010100: EEPROM_OUT = 18'b000000000000000000;
			7'b1011010: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1011011: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1011100: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1100010: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1100011: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1100100: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1101010: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1101011: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1101100: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1110010: EEPROM_OUT = 18'b000000000100000001;
			7'b1110011: EEPROM_OUT = 18'b000000000000000000;
			7'b1110100: EEPROM_OUT = 18'b000000000000000000;
			7'b1111010: EEPROM_OUT = 18'b100000000000000000;
			7'b1111011: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'b1111100: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'bxxxx101: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'bxxxx110: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;
			7'bxxxx111: EEPROM_OUT = 18'bxxxxxxxxxxxxxxxxxx;

		endcase
	end
	
endmodule